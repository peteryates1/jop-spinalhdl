--
-- bcfetch_tb.vhd
--
-- Testbench wrapper for bcfetch.vhd (bytecode fetch stage)
-- This creates a self-contained module for CocoTB testing by:
-- 1. Embedding the jbc component (bytecode RAM)
-- 2. Including the jtbl component (jump table)
-- 3. Exposing irq record fields as individual ports
-- 4. Defining required configuration constants locally
--
-- The original bcfetch.vhd depends on:
-- - jop_types.vhd (irq_bcf_type, irq_ack_type records)
-- - jop_config_global.vhd (cache configuration constants)
-- - jbc component (bytecode RAM)
-- - jtbl component (jump table - generated by Jopa)
--
-- This wrapper embeds those dependencies to simplify CocoTB testing.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bcfetch_tb is
    generic (
        jpc_width   : integer := 11;    -- address bits of java byte code pc (2KB cache)
        pc_width    : integer := 11     -- address bits of internal instruction rom
    );
    port (
        clk, reset  : in std_logic;

        -- JPC interface
        jpc_out     : out std_logic_vector(jpc_width downto 0);  -- jpc read (12-bit for 11-bit width)
        din         : in std_logic_vector(31 downto 0);          -- A from stack (for jpc_wr)
        jpc_wr      : in std_logic;                              -- write jpc from stack

        -- JBC write interface (for loading bytecode into RAM)
        bc_wr_addr  : in std_logic_vector(jpc_width-3 downto 0); -- word address
        bc_wr_data  : in std_logic_vector(31 downto 0);          -- write data (32-bit word)
        bc_wr_ena   : in std_logic;                              -- write enable

        -- Fetch control (from microcode)
        jfetch      : in std_logic;      -- fetch next bytecode
        jopdfetch   : in std_logic;      -- fetch operand byte

        -- Condition flags (from ALU/stack)
        zf, nf      : in std_logic;      -- zero flag, negative flag
        eq, lt      : in std_logic;      -- equal flag, less-than flag

        -- Branch control
        jbr         : in std_logic;      -- branch evaluation enable

        -- Interrupt interface (irq_bcf_type exposed as individual signals)
        irq_in_irq  : in std_logic;      -- interrupt request (single cycle)
        irq_in_exc  : in std_logic;      -- exception request (single cycle)
        irq_in_ena  : in std_logic;      -- global interrupt enable

        -- Interrupt acknowledge (irq_ack_type exposed as individual signals)
        irq_out_ack_irq : out std_logic; -- interrupt acknowledge
        irq_out_ack_exc : out std_logic; -- exception acknowledge

        -- Outputs
        jpaddr      : out std_logic_vector(pc_width-1 downto 0); -- microcode ROM address
        opd         : out std_logic_vector(15 downto 0);         -- operand (16-bit)

        -- Debug outputs (internal state visibility)
        dbg_jbc_data    : out std_logic_vector(7 downto 0);      -- current bytecode from RAM
        dbg_jinstr      : out std_logic_vector(7 downto 0);      -- captured instruction
        dbg_jpc_br      : out std_logic_vector(jpc_width downto 0); -- branch start PC
        dbg_jmp         : out std_logic;                         -- jump taken signal
        dbg_int_pend    : out std_logic;                         -- interrupt pending
        dbg_exc_pend    : out std_logic                          -- exception pending
    );
end bcfetch_tb;

architecture rtl of bcfetch_tb is

    --
    -- JBC component (bytecode RAM) - embedded for self-contained testbench
    -- Dual-port: 32-bit write port, 8-bit read port
    -- Registered read address, unregistered output
    --
    constant nwords : integer := 2**(jpc_width-2);
    type mem_type is array(0 to nwords-1) of std_logic_vector(31 downto 0);
    signal jbc_ram : mem_type := (others => (others => '0'));

    signal jbc_addr     : std_logic_vector(jpc_width-1 downto 0);
    signal jbc_data     : std_logic_vector(7 downto 0);
    signal jbc_addr_reg : std_logic_vector(jpc_width-1 downto 0);
    signal jbc_word     : std_logic_vector(31 downto 0);

    --
    -- Internal bcfetch signals
    --
    signal jbc_mux      : std_logic_vector(jpc_width downto 0);
    signal jbc_q        : std_logic_vector(7 downto 0);

    signal jpc          : std_logic_vector(jpc_width downto 0);
    signal jpc_br       : std_logic_vector(jpc_width downto 0);
    signal jmp_addr     : std_logic_vector(jpc_width downto 0);

    signal jinstr       : std_logic_vector(7 downto 0);
    signal tp           : std_logic_vector(3 downto 0);
    signal jmp          : std_logic;

    signal jopd         : std_logic_vector(15 downto 0);

    -- Interrupt handling signals
    signal int_pend     : std_logic;
    signal int_req      : std_logic;
    signal int_taken    : std_logic;

    signal exc_pend     : std_logic;
    signal exc_taken    : std_logic;

    signal bytecode     : std_logic_vector(7 downto 0);

    -- Jump table output
    signal jtbl_addr    : std_logic_vector(pc_width-1 downto 0);

begin

    --
    -- JBC RAM implementation (embedded)
    -- Write: 32-bit words at word address
    -- Read: 8-bit bytes at byte address (registered address, unregistered output)
    --
    process(clk)
    begin
        if rising_edge(clk) then
            -- Write port (32-bit)
            if bc_wr_ena = '1' then
                jbc_ram(to_integer(unsigned(bc_wr_addr))) <= bc_wr_data;
            end if;

            -- Register read address
            jbc_addr_reg <= jbc_addr;
        end if;
    end process;

    -- Read port - word lookup
    jbc_word <= jbc_ram(to_integer(unsigned(jbc_addr_reg(jpc_width-1 downto 2))));

    -- Byte selection mux (unregistered output)
    process(jbc_addr_reg, jbc_word)
    begin
        case jbc_addr_reg(1 downto 0) is
            when "11" =>
                jbc_data <= jbc_word(31 downto 24);
            when "10" =>
                jbc_data <= jbc_word(23 downto 16);
            when "01" =>
                jbc_data <= jbc_word(15 downto 8);
            when "00" =>
                jbc_data <= jbc_word(7 downto 0);
            when others =>
                jbc_data <= (others => '0');
        end case;
    end process;

    --
    -- Jump table (jtbl) - instantiate generated component
    --
    jt: entity work.jtbl
        port map (
            bcode    => bytecode,
            int_pend => int_req,
            exc_pend => exc_pend,
            q        => jtbl_addr
        );

    --
    -- Interrupt processing
    --
    process(clk, reset)
    begin
        if (reset = '1') then
            int_pend <= '0';
            exc_pend <= '0';
        elsif rising_edge(clk) then
            if irq_in_irq = '1' then
                int_pend <= '1';
            elsif int_taken = '1' then
                int_pend <= '0';
            end if;

            if irq_in_exc = '1' then
                exc_pend <= '1';
            elsif exc_taken = '1' then
                exc_pend <= '0';
            end if;
        end if;
    end process;

    int_req <= int_pend and irq_in_ena;
    int_taken <= int_req and jfetch;
    exc_taken <= exc_pend and jfetch;

    irq_out_ack_irq <= int_taken;
    irq_out_ack_exc <= exc_taken;

    --
    -- Bytecode to jump table
    --
    bytecode <= jbc_q;
    jpaddr <= jtbl_addr;

    jbc_addr <= jbc_mux(jpc_width-1 downto 0);
    jbc_q <= jbc_data;

    --
    -- Branch type decode (registered)
    --
    process(clk, jinstr)
    begin
        if rising_edge(clk) then
            case jinstr is
                when "10100101" => tp <= "1111";    -- if_acmpeq
                when "10100110" => tp <= "0000";    -- if_acmpne
                when "11000110" => tp <= "1001";    -- ifnull
                when "11000111" => tp <= "1010";    -- ifnonnull
                when others => tp <= jinstr(3 downto 0);
            end case;
        end if;
    end process;

    --
    -- Branch condition evaluation (combinational)
    --
    process(tp, jbr, zf, nf, eq, lt)
    begin
        jmp <= '0';
        if (jbr = '1') then
            case tp is
                when "1001" =>          -- ifeq, ifnull
                    if (zf = '1') then
                        jmp <= '1';
                    end if;
                when "1010" =>          -- ifne, ifnonnull
                    if (zf = '0') then
                        jmp <= '1';
                    end if;
                when "1011" =>          -- iflt
                    if (nf = '1') then
                        jmp <= '1';
                    end if;
                when "1100" =>          -- ifge
                    if (nf = '0') then
                        jmp <= '1';
                    end if;
                when "1101" =>          -- ifgt
                    if (zf = '0' and nf = '0') then
                        jmp <= '1';
                    end if;
                when "1110" =>          -- ifle
                    if (zf = '1' or nf = '1') then
                        jmp <= '1';
                    end if;
                when "1111" =>          -- if_icmpeq, if_acmpeq
                    if (eq = '1') then
                        jmp <= '1';
                    end if;
                when "0000" =>          -- if_icmpne, if_acmpne
                    if (eq = '0') then
                        jmp <= '1';
                    end if;
                when "0001" =>          -- if_icmplt
                    if (lt = '1') then
                        jmp <= '1';
                    end if;
                when "0010" =>          -- if_icmpge
                    if (lt = '0') then
                        jmp <= '1';
                    end if;
                when "0011" =>          -- if_icmpgt
                    if (eq = '0' and lt = '0') then
                        jmp <= '1';
                    end if;
                when "0100" =>          -- if_icmple
                    if (eq = '1' or lt = '1') then
                        jmp <= '1';
                    end if;
                when "0111" =>          -- goto
                    jmp <= '1';
                when others =>
                    null;
            end case;
        end if;
    end process;

    --
    -- JBC read address mux
    --
    process(din, jpc, jmp_addr, jopd, jfetch, jopdfetch, jmp)
    begin
        if (jmp = '1') then
            jbc_mux <= jmp_addr;
        elsif (jfetch = '1' or jopdfetch = '1') then
            jbc_mux <= std_logic_vector(unsigned(jpc) + 1);
        else
            jbc_mux <= jpc;
        end if;
    end process;

    --
    -- JPC update logic
    --
    process(clk, reset)
    begin
        if (reset = '1') then
            jpc <= std_logic_vector(to_unsigned(0, jpc_width+1));
        elsif rising_edge(clk) then
            if (jpc_wr = '1') then
                jpc <= din(jpc_width downto 0);
            elsif (jmp = '1') then
                jpc <= jmp_addr;
            elsif (jfetch = '1' or jopdfetch = '1') then
                jpc <= std_logic_vector(unsigned(jpc) + 1);
            else
                jpc <= jpc;
            end if;
        end if;
    end process;

    jpc_out <= jpc;

    --
    -- Branch address calculation and instruction capture
    --
    process(clk)
        variable branch_offset : std_logic_vector(jpc_width downto 0);
    begin
        if rising_edge(clk) then
            -- Branch target: jpc_br + signed(jopd_high & jbc_q)
            -- Build the offset by concatenating operand high bits with current bytecode
            branch_offset := jopd(jpc_width-8 downto 0) & jbc_q;
            jmp_addr <= std_logic_vector(unsigned(jpc_br) + unsigned(branch_offset));

            if (jfetch = '1') then
                jpc_br <= jpc;          -- save start address for branch
                jinstr <= jbc_q;        -- capture bytecode
            end if;
        end if;
    end process;

    --
    -- Operand accumulation
    --
    process(clk, reset)
    begin
        if (reset = '1') then
            jopd <= (others => '0');
        elsif rising_edge(clk) then
            jopd(7 downto 0) <= jbc_q;  -- low byte always updates
            if (jopdfetch = '1') then
                jopd(15 downto 8) <= jopd(7 downto 0);  -- shift low to high
            end if;
        end if;
    end process;

    opd <= jopd;

    --
    -- Debug outputs
    --
    dbg_jbc_data <= jbc_q;
    dbg_jinstr <= jinstr;
    dbg_jpc_br <= jpc_br;
    dbg_jmp <= jmp;
    dbg_int_pend <= int_pend;
    dbg_exc_pend <= exc_pend;

end rtl;
