`timescale 1ns/1ps

module tb_jop_gc_sdram;

  // Clock and reset
  reg clk = 0;
  reg reset = 1;

  // 100 MHz clock (10ns period)
  always #5 clk = ~clk;

  // Reset sequence: hold reset for 100ns then release
  initial begin
    reset = 1;
    #100;
    reset = 0;
  end

  // DUT outputs
  wire [10:0] pc;
  wire [11:0] jpc;
  wire [9:0]  instr;
  wire        jfetch;
  wire        jopdfetch;
  wire [31:0] aout;
  wire [31:0] bout;
  wire        memBusy;
  wire [7:0]  uartTxData;
  wire        uartTxValid;
  wire        ioWr;
  wire [7:0]  ioAddr;
  wire [31:0] ioWrData;

  // BMB debug
  wire        bmbCmdValid;
  wire        bmbCmdReady;
  wire [25:0] bmbCmdAddr;
  wire [0:0]  bmbCmdOpcode;
  wire        bmbRspValid;
  wire [31:0] bmbRspData;

  // SDRAM interface (directly wired between DUT and SDRAM model)
  wire [12:0] sdram_addr;
  wire [1:0]  sdram_ba;
  wire        sdram_casn;
  wire        sdram_cke;
  wire        sdram_csn;
  wire [15:0] sdram_dq;
  wire [1:0]  sdram_dqm;
  wire        sdram_rasn;
  wire        sdram_wen;

  // Instantiate DUT
  JopCoreWithSdramTestHarness dut (
    .clk                (clk),
    .reset              (reset),
    .io_sdram_ADDR      (sdram_addr),
    .io_sdram_BA        (sdram_ba),
    .io_sdram_CASn      (sdram_casn),
    .io_sdram_CKE       (sdram_cke),
    .io_sdram_CSn       (sdram_csn),
    .io_sdram_DQ        (sdram_dq),
    .io_sdram_DQM       (sdram_dqm),
    .io_sdram_RASn      (sdram_rasn),
    .io_sdram_WEn       (sdram_wen),
    .io_pc              (pc),
    .io_jpc             (jpc),
    .io_instr           (instr),
    .io_jfetch          (jfetch),
    .io_jopdfetch       (jopdfetch),
    .io_aout            (aout),
    .io_bout            (bout),
    .io_memBusy         (memBusy),
    .io_uartTxData      (uartTxData),
    .io_uartTxValid     (uartTxValid),
    .io_ioWr            (ioWr),
    .io_ioAddr          (ioAddr),
    .io_ioWrData        (ioWrData),
    .io_bmbCmdValid     (bmbCmdValid),
    .io_bmbCmdReady     (bmbCmdReady),
    .io_bmbCmdAddr      (bmbCmdAddr),
    .io_bmbCmdOpcode    (bmbCmdOpcode),
    .io_bmbRspValid     (bmbRspValid),
    .io_bmbRspData      (bmbRspData)
  );

  // Instantiate SDRAM model with timing assertions
  // W9825G6JH6 parameters: 13-bit row, 9-bit col, CAS=3, 8MB
  sdram_model #(
    .ROW_BITS   (13),
    .COL_BITS   (9),
    .BANK_BITS  (2),
    .DQ_BITS    (16),
    .CAS        (3),
    .tRP_CYC    (2),    // 20ns / 10ns = 2 cycles
    .tRCD_CYC   (2),    // 20ns / 10ns = 2 cycles
    .tRAS_CYC   (5),    // 45ns / 10ns = 4.5, round up = 5
    .tRC_CYC    (6),    // 65ns / 10ns = 6.5, round up = 7 but SdramCtrl uses 6
    .tWR_CYC    (1),    // 1 cycle write recovery (tDPL)
    .tRFC_CYC   (6),    // 66ns / 10ns = 6.6, round up = 7 but use 6
    .MEM_BYTES  (8*1024*1024)  // 8MB (W9825G6JH6 = 256Mbit / 8 / 2 chips? = 8MB per chip actually 32MB but we use 8MB for the model)
  ) sdram (
    .clk    (clk),
    .cke    (sdram_cke),
    .cs_n   (sdram_csn),
    .ras_n  (sdram_rasn),
    .cas_n  (sdram_casn),
    .we_n   (sdram_wen),
    .ba     (sdram_ba),
    .addr   (sdram_addr),
    .dqm    (sdram_dqm),
    .dq     (sdram_dq)
  );

  // Load SDRAM with program data
  // The sdram_init.hex file is generated by JopSmallGcSdramQuestaGen
  // It contains 32-bit words; we need to convert to the SDRAM model's byte-addressed memory
  reg [31:0] init_data [0:32767];  // 128KB / 4 = 32K words
  integer init_i;

  initial begin
    $readmemh("sdram_init.hex", init_data);
    // Convert 32-bit words to byte-addressed SDRAM memory
    // SDRAM model address mapping: {row, bank, column} * 2 bytes
    // But for initialization, we use linear byte addressing
    for (init_i = 0; init_i < 32768; init_i = init_i + 1) begin
      // Little-endian byte order (matching SpinalHDL SdramModel)
      sdram.mem[init_i*4 + 0] = init_data[init_i][7:0];
      sdram.mem[init_i*4 + 1] = init_data[init_i][15:8];
      sdram.mem[init_i*4 + 2] = init_data[init_i][23:16];
      sdram.mem[init_i*4 + 3] = init_data[init_i][31:24];
    end
    $display("SDRAM initialized: 32768 words from sdram_init.hex");
    // Verify initialization
    $display("  init_data[0] = %h (expect 00002065)", init_data[0]);
    $display("  init_data[1] = %h (expect 0000144f)", init_data[1]);
    $display("  sdram.mem[0:3] = %h %h %h %h (expect 65 20 00 00)",
             sdram.mem[0], sdram.mem[1], sdram.mem[2], sdram.mem[3]);
    $display("  sdram.mem[4:7] = %h %h %h %h (expect 4f 14 00 00)",
             sdram.mem[4], sdram.mem[5], sdram.mem[6], sdram.mem[7]);
  end

  // Cycle counter
  integer cycle_count = 0;
  integer max_cycles = 20000000;  // 20M cycles

  // UART tracking
  integer found_gc_start = 0;
  integer found_r14 = 0;
  integer extra_cycles = 0;

  // BMB transaction monitoring
  integer bmb_reads = 0;
  integer bmb_writes = 0;
  integer bmb_stalls = 0;  // cycles where cmd.valid && !cmd.ready

  // Main simulation loop
  always @(posedge clk) begin
    if (!reset) begin
      cycle_count <= cycle_count + 1;

      // Monitor UART output
      if (uartTxValid) begin
        if (uartTxData >= 32 && uartTxData < 127)
          $write("%c", uartTxData);
        else if (uartTxData == 8'h0A)
          $write("\n");
        else if (uartTxData == 8'h0D)
          ; // skip CR
        else
          $write(".");
      end

      // Monitor BMB transactions (detailed logging for first 50 transactions)
      if (bmbCmdValid && bmbCmdReady) begin
        if (bmbCmdOpcode == 0) begin
          bmb_reads <= bmb_reads + 1;
          if (bmb_reads < 50)
            $display("[%0d] BMB READ  addr=%h", cycle_count, bmbCmdAddr);
        end else begin
          bmb_writes <= bmb_writes + 1;
          if (bmb_writes < 50)
            $display("[%0d] BMB WRITE addr=%h", cycle_count, bmbCmdAddr);
        end
      end
      if (bmbCmdValid && !bmbCmdReady) begin
        bmb_stalls <= bmb_stalls + 1;
      end

      // Monitor BMB responses
      if (bmbRspValid && (bmb_reads + bmb_writes < 55)) begin
        $display("[%0d] BMB RSP   data=%h", cycle_count, bmbRspData);
      end

      // Monitor SDRAM DQ bus and control signals around init
      if (cycle_count > 32825 && cycle_count < 32850) begin
        $display("[%0d] SDRAM csn=%b rasn=%b casn=%b wen=%b ba=%b addr=%h dq=%h dqm=%b model_oe=%b model_drive=%h pipe_v2=%b pipe_d2=%h dut_dq_we0=%b",
                 cycle_count, sdram_csn, sdram_rasn, sdram_casn, sdram_wen,
                 sdram_ba, sdram_addr, sdram_dq, sdram_dqm,
                 sdram.dq_oe_neg, sdram.dq_drive,
                 sdram.read_pipe_valid[2], sdram.read_pipe_data[2],
                 dut._zz_io_sdram_DQ);
      end

      // Progress report every 100k cycles
      if (cycle_count > 0 && cycle_count % 100000 == 0) begin
        $display("\n[%0d] PC=%h JPC=%h memBusy=%b reads=%0d writes=%0d stalls=%0d violations=%0d",
                 cycle_count, pc, jpc, memBusy,
                 bmb_reads, bmb_writes, bmb_stalls,
                 sdram.timing_violations);
      end

      // Timeout
      if (cycle_count >= max_cycles) begin
        $display("\n\n=== TIMEOUT after %0d cycles ===", cycle_count);
        $display("BMB: %0d reads, %0d writes, %0d stall cycles", bmb_reads, bmb_writes, bmb_stalls);
        $display("SDRAM: %0d timing violations", sdram.timing_violations);
        $display("SDRAM: %0d activates, %0d precharges, %0d refreshes",
                 sdram.total_activates, sdram.total_precharges, sdram.total_refreshes);
        if (sdram.timing_violations > 0)
          $display("*** TIMING VIOLATIONS DETECTED — check log above ***");
        else
          $display("No SDRAM timing violations detected.");
        $finish;
      end
    end
  end

endmodule
